module Lab1 (
    input butnS2_n,
    output led
);

assign led = butnS2_n;

endmodule
